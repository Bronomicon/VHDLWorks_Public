ENTITY TB_AW IS

END TB_AW;


ARCHITECTURE AW_BEH OF TB_AW IS
	
	COMPONENT AW IS
	GENERIC	(N: Integer:=4); --Bitmenge des Addierwerkes
	PORT		(NumberA:	IN BIT_VECTOR (N-1 DOWNTO 0);
				 NumberB:	IN BIT_VECTOR (N-1 DOWNTO 0);
				 NumberC:	OUT BIT_VECTOR (N DOWNTO 0));
	END COMPONENT;
	
	
   SIGNAL NumberA_test: BIT_VECTOR (3 DOWNTO 0);
	SIGNAL NumberB_test: BIT_VECTOR (3 DOWNTO 0);
	SIGNAL NumberC_test: BIT_VECTOR (4 DOWNTO 0);

	
	BEGIN
	AW_TEST: AW PORT MAP(NumberA_test, NumberB_test, NumberC_test);
	
	NumberA_test <= "0000", "0001" AFTER 10ns, "1011" AFTER 20ns, "1111" AFTER 30ns;
	NumberB_test <= "0000", "0001" AFTER 10ns, "1011" AFTER 20ns, "1111" AFTER 30ns;

END AW_BEH;
		
		